--							dcdr01.vhd
-- Декодер-формирователь управляющих данных для конечного автомата,
-- выдающего на светодиод серию из пяти вспышек, соответствующих
-- пятибитному двоичному числу (используется для идентификации версии
-- прошивки ПЛИС).

-- Разработан для проекта преобразователя интерфейса ISDN-IP 06.11.2023

entity dcdr01 is
port(
-- CIN[4..0] - Пятибитное двоичное число, отображаемое на одиночном
-- светодиоде в виде последовательности вспышек длительностью 0,25 с
-- (логический 0) и 0,75 с (логическая 1), разделенных интервалами
-- по 0,5 с. Для работы логической схемы является задаваемой
-- пользователем константой
--
-- ST[2..0] - Трехбитное двоичное число, обозначающее номер генерируемой
-- вспышки в последовательности
--
-- V0_EQU[4..0] - Пятибитное двоичное число, обозначающее номер такта,
-- на котором происходит переключение выдаваемого сигнала в логический 0
--
-- V1_EQU[4..0] - Пятибитное двоичное число, обозначающее номер такта,
-- на котором происходит переключение выдаваемого сигнала в логическую 1
--
-- NULL_EQU[4..0] - - Пятибитное двоичное число, обозначающее номер
-- такта, на котором происходит установка счетчика-формирователя
-- в нулевое состояние

CIN: in bit_vector (4 downto 0);
ST: in bit_vector (2 downto 0);
V0_EQU: out bit_vector (4 downto 0);
V1_EQU: out bit_vector (4 downto 0);
NULL_EQU: out bit_vector (4 downto 0)
); -- port
end dcdr01;

architecture ttable of dcdr01 is
	signal TMP_IN: bit_vector(7 downto 0);
	signal TMP_OUT: bit_vector(14 downto 0);

-- Лог.0 (NULL_EQU = 5 b'00101') (V0_EQU = 3 b'00011') (V1_EQU = 1 b'00001')
--
--				Значение счетчика, при котором происходит
-- 				переключение в логический 0			  │						  ┐
--													  │
--				Значение счетчика,					  │
--				при котором происходит сброс в 0 ┐	  │
--											   ┌─┴─┐┌─┴─┐┌─┴─┐
	constant LOG_0: bit_vector(14 downto 0) :="001010001100001";
	
-- Лог.1 (NULL_EQU = 9 b'01001') (V0_EQU = 7 b'00111') (V1_EQU = 1 b'00001')	
	constant LOG_1: bit_vector(14 downto 0) :="010010011100001";
	
begin

-- Объединяем в одном векторе входные (ST с CIN) и выходные (V1_EQU,
-- V0_EQU, NULL_EQU) битовые векторы для использования оператором
-- select. При анализе/корректировке кода ОСОБОЕ ВНИМАНИЕ ОБРАТИТЬ
-- на последовательность битов и переменных в объединенных векторах.

-- Входы
	TMP_IN(7 downto 3) <= CIN;
	TMP_IN(2 downto 0) <= ST;
	
-- Выходы	
	NULL_EQU(4 downto 0) <= TMP_OUT(14 downto 10);
	V0_EQU(4 downto 0) <= TMP_OUT(9 downto 5);
	V1_EQU(4 downto 0) <= TMP_OUT(4 downto 0);

-- Определяем таблицу истинности
	with TMP_IN select TMP_OUT <=

--	   TMP_OUT		 TMP_IN
-- 0 b'00000'
--	 				  ┌───── Кодируемое последовательностью число 
--					  │	  ┌─ Номер вспышки
--					┌─┴─┐┌┴┐
		LOG_0 when "00000000", -- 0 MSB выдается первым
		LOG_0 when "00000001", -- 0
		LOG_0 when "00000010", -- 0
		LOG_0 when "00000011", -- 0
		LOG_0 when "00000100", -- 0 LSB выдается последним
-- 1 b'00001'
		LOG_0 when "00001000", -- 0 MSB выдается первым
		LOG_0 when "00001001", -- 0
		LOG_0 when "00001010", -- 0
		LOG_0 when "00001011", -- 0
		LOG_1 when "00001100", -- 1 LSB выдается последним
-- 2 b'00010'
		LOG_0 when "00010000", -- 0 MSB выдается первым
		LOG_0 when "00010001", -- 0
		LOG_0 when "00010010", -- 0
		LOG_1 when "00010011", -- 1
		LOG_0 when "00010100", -- 0 LSB выдается последним
-- 3 b'00011'
		LOG_0 when "00011000", -- 0 MSB выдается первым
		LOG_0 when "00011001", -- 0
		LOG_0 when "00011010", -- 0
		LOG_1 when "00011011", -- 1
		LOG_1 when "00011100", -- 1 LSB выдается последним
-- 4 b'00100'
		LOG_0 when "00100000", -- 0 MSB выдается первым
		LOG_0 when "00100001", -- 0
		LOG_1 when "00100010", -- 1
		LOG_0 when "00100011", -- 0
		LOG_0 when "00100100", -- 0 LSB выдается последним
-- 5 b'00101'
		LOG_0 when "00101000", -- 0 MSB выдается первым
		LOG_0 when "00101001", -- 0
		LOG_1 when "00101010", -- 1
		LOG_0 when "00101011", -- 0
		LOG_1 when "00101100", -- 1 LSB выдается последним
-- 6 b'00110'
		LOG_0 when "00110000", -- 0 MSB выдается первым
		LOG_0 when "00110001", -- 0
		LOG_1 when "00110010", -- 1
		LOG_1 when "00110011", -- 1
		LOG_0 when "00110100", -- 0 LSB выдается последним
-- 7 b'00111'
		LOG_0 when "00111000", -- 0 MSB выдается первым
		LOG_0 when "00111001", -- 0
		LOG_1 when "00111010", -- 1
		LOG_1 when "00111011", -- 1
		LOG_1 when "00111100", -- 1 LSB выдается последним
-- 8 b'01000'
		LOG_0 when "01000000", -- 0 MSB выдается первым
		LOG_1 when "01000001", -- 1
		LOG_0 when "01000010", -- 0
		LOG_0 when "01000011", -- 0
		LOG_0 when "01000100", -- 0 LSB выдается последним
-- 9 b'01001'
		LOG_0 when "01001000", -- 0 MSB выдается первым
		LOG_1 when "01001001", -- 1
		LOG_0 when "01001010", -- 0
		LOG_0 when "01001011", -- 0
		LOG_1 when "01001100", -- 1 LSB выдается последним
-- 10 b'01010'
		LOG_0 when "01010000", -- 0 MSB выдается первым
		LOG_1 when "01010001", -- 1
		LOG_0 when "01010010", -- 0
		LOG_1 when "01010011", -- 1
		LOG_0 when "01010100", -- 0 LSB выдается последним
-- 11 b'01011'
		LOG_0 when "01011000", -- 0 MSB выдается первым
		LOG_1 when "01011001", -- 1
		LOG_0 when "01011010", -- 0
		LOG_1 when "01011011", -- 1
		LOG_1 when "01011100", -- 1 LSB выдается последним
-- 12 b'01100'
		LOG_0 when "01100000", -- 0 MSB выдается первым
		LOG_1 when "01100001", -- 1
		LOG_1 when "01100010", -- 1
		LOG_0 when "01100011", -- 0
		LOG_0 when "01100100", -- 0 LSB выдается последним
-- 13 b'01101'
		LOG_0 when "01101000", -- 0 MSB выдается первым
		LOG_1 when "01101001", -- 1
		LOG_1 when "01101010", -- 1
		LOG_0 when "01101011", -- 0
		LOG_1 when "01101100", -- 1 LSB выдается последним
-- 14 b'01110'
		LOG_0 when "01110000", -- 0 MSB выдается первым
		LOG_1 when "01110001", -- 1
		LOG_1 when "01110010", -- 1
		LOG_1 when "01110011", -- 1
		LOG_0 when "01110100", -- 0 LSB выдается последним
-- 15 b'01111'
		LOG_0 when "01111000", -- 0 MSB выдается первым
		LOG_1 when "01111001", -- 1
		LOG_1 when "01111010", -- 1
		LOG_1 when "01111011", -- 1
		LOG_1 when "01111100", -- 1 LSB выдается последним
-- 16 b'10000'
		LOG_1 when "10000000", -- 1 MSB выдается первым
		LOG_0 when "10000001", -- 0
		LOG_0 when "10000010", -- 0
		LOG_0 when "10000011", -- 0
		LOG_0 when "10000100", -- 0 LSB выдается последним
-- 17 b'10001'
		LOG_1 when "10001000", -- 1 MSB выдается первым
		LOG_0 when "10001001", -- 0
		LOG_0 when "10001010", -- 0
		LOG_0 when "10001011", -- 0
		LOG_1 when "10001100", -- 1 LSB выдается последним
-- 18 b'10010'
		LOG_1 when "10010000", -- 1 MSB выдается первым
		LOG_0 when "10010001", -- 0
		LOG_0 when "10010010", -- 0
		LOG_1 when "10010011", -- 1
		LOG_0 when "10010100", -- 0 LSB выдается последним
-- 19 b'10011'
		LOG_1 when "10011000", -- 1 MSB выдается первым
		LOG_0 when "10011001", -- 0
		LOG_0 when "10011010", -- 0
		LOG_1 when "10011011", -- 1
		LOG_1 when "10011100", -- 1 LSB выдается последним
-- 20 b'00100'
		LOG_1 when "10100000", -- 1 MSB выдается первым
		LOG_0 when "10100001", -- 0
		LOG_1 when "10100010", -- 1
		LOG_0 when "10100011", -- 0
		LOG_0 when "10100100", -- 0 LSB выдается последним
-- 21 b'00101'
		LOG_1 when "10101000", -- 1 MSB выдается первым
		LOG_0 when "10101001", -- 0
		LOG_1 when "10101010", -- 1
		LOG_0 when "10101011", -- 0
		LOG_1 when "10101100", -- 1 LSB выдается последним
-- 22 b'00110'
		LOG_1 when "10110000", -- 1 MSB выдается первым
		LOG_0 when "10110001", -- 0
		LOG_1 when "10110010", -- 1
		LOG_1 when "10110011", -- 1
		LOG_0 when "10110100", -- 0 LSB выдается последним
-- 23 b'00111'
		LOG_1 when "10111000", -- 1 MSB выдается первым
		LOG_0 when "10111001", -- 0
		LOG_1 when "10111010", -- 1
		LOG_1 when "10111011", -- 1
		LOG_1 when "10111100", -- 1 LSB выдается последним
-- 24 b'01000'
		LOG_1 when "11000000", -- 1 MSB выдается первым
		LOG_1 when "11000001", -- 1
		LOG_0 when "11000010", -- 0
		LOG_0 when "11000011", -- 0
		LOG_0 when "11000100", -- 0 LSB выдается последним
-- 25 b'01001'
		LOG_1 when "11001000", -- 1 MSB выдается первым
		LOG_1 when "11001001", -- 1
		LOG_0 when "11001010", -- 0
		LOG_0 when "11001011", -- 0
		LOG_1 when "11001100", -- 1 LSB выдается последним
-- 26 b'01010'
		LOG_1 when "11010000", -- 1 MSB выдается первым
		LOG_1 when "11010001", -- 1
		LOG_0 when "11010010", -- 0
		LOG_1 when "11010011", -- 1
		LOG_0 when "11010100", -- 0 LSB выдается последним
-- 27 b'01011'
		LOG_1 when "11011000", -- 1 MSB выдается первым
		LOG_1 when "11011001", -- 1
		LOG_0 when "11011010", -- 0
		LOG_1 when "11011011", -- 1
		LOG_1 when "11011100", -- 1 LSB выдается последним
-- 28 b'01100'
		LOG_1 when "11100000", -- 1 MSB выдается первым
		LOG_1 when "11100001", -- 1
		LOG_1 when "11100010", -- 1
		LOG_0 when "11100011", -- 0
		LOG_0 when "11100100", -- 0 LSB выдается последним
-- 29 b'01101'
		LOG_1 when "11101000", -- 1 MSB выдается первым
		LOG_1 when "11101001", -- 1
		LOG_1 when "11101010", -- 1
		LOG_0 when "11101011", -- 0
		LOG_1 when "11101100", -- 1 LSB выдается последним
-- 30 b'01110'
		LOG_1 when "11110000", -- 1 MSB выдается первым
		LOG_1 when "11110001", -- 1
		LOG_1 when "11110010", -- 1
		LOG_1 when "11110011", -- 1
		LOG_0 when "11110100", -- 0 LSB выдается последним
-- 31 b'01111'
		LOG_1 when "11111000", -- 1 MSB выдается первым
		LOG_1 when "11111001", -- 1
		LOG_1 when "11111010", -- 1
		LOG_1 when "11111011", -- 1
		LOG_1 when "11111100", -- 1 LSB выдается последним

		"111111111111111" when others;
end ttable;
