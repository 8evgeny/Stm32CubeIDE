DCE01_SFL_inst : DCE01_SFL PORT MAP (
		noe_in	 => noe_in_sig
	);
